interface intf1(input logic clk);
logic signed [4:0] A;
logic signed [4:0] B;
logic signed [2:0] a_op;
logic signed [1:0] b_op;
logic a_en;
logic b_en;
logic ALU_en;
logic rst_n;
logic signed [5:0] C;

endinterface